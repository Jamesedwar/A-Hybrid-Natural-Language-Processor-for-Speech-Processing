module word_Library(clock, enable, address, out);
input          clock;
input         enable;
input   [7:0]address;
output     [79:0]out;

reg [79:0]mem[0:255];
reg        [79:0]out;
always@(posedge clock or negedge enable)
begin
if(enable == 0)
begin
out<=80'd0;
mem[0]<=80'h00000000000000000020;
//1st Sentence
mem[1]<=80'h00000053616d73756e67;
mem[2]<=80'h00000000000000006973;
mem[3]<=80'h0000006c6f6361746564;
mem[4]<=80'h0000000000000000696e;
mem[5]<=80'h0000000000536f757468;
mem[6]<=80'h00000000004b6f726561;
mem[7]<=80'h0000000000000000002e;
mem[8]<=80'h00000000005768657265;
mem[9]<=80'h00000000000000006973;
mem[10]<=80'h00000053616d73756e67;
mem[11]<=80'h0000006c6f6361746564;
mem[12]<=80'h0000000000000000003f;
//2nd Sentence
mem[13]<=80'h000000000000004c6565;
mem[14]<=80'h00000000004279756e67;
mem[15]<=80'h00000000000000006973;
mem[16]<=80'h00000000000000746865;
mem[17]<=80'h000000666f756e646572;
mem[18]<=80'h00000000000000006f66;
mem[19]<=80'h00000053616d73756e67;
mem[20]<=80'h0000000000000000002e;
mem[21]<=80'h0000000000000057686f;
mem[22]<=80'h00000000000000006973;
mem[23]<=80'h00000000000000746865;
mem[24]<=80'h000000666f756e646572;
mem[25]<=80'h00000000000000006f66;
mem[26]<=80'h00000053616d73756e67;
mem[27]<=80'h0000000000000000003f;
//3rd Sentence
mem[28]<=80'h00000000000000546865;
mem[29]<=80'h00000063757272656e74;
mem[30]<=80'h0000000000666f637573;
mem[31]<=80'h00000000000000006f66;
mem[32]<=80'h00000053616d73756e67;
mem[33]<=80'h00000000000000006973;
mem[34]<=80'h0000000000536d617274;
mem[35]<=80'h0000000070686f6e6573;
mem[36]<=80'h0000000000000000002e;
mem[37]<=80'h00000000000057686174;
mem[38]<=80'h00000000000000006973;
mem[39]<=80'h00000000000000546865;
mem[40]<=80'h0000000000666f637573;
mem[41]<=80'h00000000000000006f66;
mem[42]<=80'h00000053616d73756e67;
mem[43]<=80'h0000000000000000003f;

//4th Sentence
mem[44]<=80'h00000000000000005336;
mem[45]<=80'h00000000000000776173;
mem[46]<=80'h000072656c6561736564;
mem[47]<=80'h0000000000000000696e;
mem[48]<=80'h00000000000032303135;
mem[49]<=80'h0000000000000000002e;
mem[50]<=80'h0000000000005768656e;
mem[51]<=80'h00000000000000776173;
mem[52]<=80'h00000000000000005336;
mem[53]<=80'h000072656c6561736564;
mem[54]<=80'h0000000000000000003f;

// 5th Sentence
mem[55]<=80'h00000000000000005336;
mem[56]<=80'h00000000000000686173;
mem[57]<=80'h000000416e64726f6964;
mem[58]<=80'h00000000000000004f53;
mem[59]<=80'h0000000000000000002e;
mem[60]<=80'h00000000005768696368;
mem[61]<=80'h00000000000000004f53;
mem[62]<=80'h00000000000000006973;
mem[63]<=80'h00000070726573656e74;
mem[64]<=80'h0000000000000000696e;
mem[65]<=80'h00000000000000005336;
mem[66]<=80'h0000000000000000003f;


//6th Sentence
mem[67]<=80'h00000053616d73756e67;
mem[68]<=80'h00000000000000006973;
mem[69]<=80'h00000000000000000061;
mem[70]<=80'h00000000676c6f62616c;
mem[71]<=80'h000000636f6d70616e79;
mem[72]<=80'h0000000000000000002e;
mem[73]<=80'h00000000000000004973;
mem[74]<=80'h00000053616d73756e67;
mem[75]<=80'h00000000000000000061;
mem[76]<=80'h00006e6174696f6e616c;
mem[77]<=80'h000000636f6d70616e79;
mem[78]<=80'h0000000000000000003f;

//7th Sentence
mem[79]<=80'h0000000000004d61696e;
mem[80]<=80'h636f6d70657469746f72;
mem[81]<=80'h00000000000000006f66;
mem[82]<=80'h00000053616d73756e67;
mem[83]<=80'h00000000000000006973;
mem[84]<=80'h00000000004170706c65;
mem[85]<=80'h0000000000000000002e;
mem[86]<=80'h00000000000000546865;
mem[87]<=80'h0000000000004d61696e;
mem[88]<=80'h636f6d70657469746f72;  
mem[89]<=80'h00000000000000006f66;   
mem[90]<=80'h00000053616d73756e67;
mem[91]<=80'h0000000000000000003f;

//8th Sentence
mem[92]<=80'h00000000000000005336;
mem[93]<=80'h0000000000636f737473;
mem[94]<=80'h00000000000031303030;
mem[95]<=80'h000052696e6767697473;
mem[96]<=80'h0000000000000000002e;
mem[97]<=80'h00000000000000486f77;
mem[98]<=80'h0000000000006d756368;
mem[99]<=80'h000000000000646f6573;
mem[100]<=80'h00000000000000005336;
mem[101]<=80'h000000000000636f7374;
mem[102]<=80'h0000000000000000003f;

//9th Sentence
mem[103]<=80'h00000000000000005336;
mem[104]<=80'h0000000000000052414d;
mem[105]<=80'h00000000000073697a65;
mem[106]<=80'h00000000000000006973;
mem[107]<=80'h00000000000000000033;
mem[108]<=80'h00000000000000004742;
mem[109]<=80'h0000000000000000002e;
mem[110]<=80'h00000000000054656c6c;
mem[111]<=80'h00000000000000746865;
mem[112]<=80'h0000000000000052414d;
mem[113]<=80'h00000000000073697a65;
mem[114]<=80'h00000000000000006f66;
mem[115]<=80'h00000000000000005336;
mem[116]<=80'h0000000000000000003f;

//10th Sentence
mem[117]<=80'h00000041697261736961;
mem[118]<=80'h0000000000006d61696e;
mem[119]<=80'h000000006f6666696365;
mem[120]<=80'h00000000000000006973;
mem[121]<=80'h0000006c6f6361746564;
mem[122]<=80'h0000000000000000696e;
mem[123]<=80'h00000000537562616e67;
mem[124]<=80'h0000000000004a617961;
mem[125]<=80'h0000000000000000002e;
mem[126]<=80'h00004169726173696173;
mem[127]<=80'h0000000000006d61696e;
mem[128]<=80'h000000006f6666696365;
mem[129]<=80'h00000000000000006973;
mem[130]<=80'h0000006c6f6361746564;
mem[131]<=80'h0000000000000000696e;
mem[132]<=80'h0000000000000000003f;

//11th Sentence
mem[133]<=80'h0000000000414b303231;
mem[134]<=80'h00000061727269766573;
mem[135]<=80'h0000000000000000696e;
mem[136]<=80'h00000000000000000034;
mem[137]<=80'h0000000000686f757273;
mem[138]<=80'h0000000000000000002e;
mem[139]<=80'h000000414b3032312773;
mem[140]<=80'h0000006172726976616c;
mem[141]<=80'h00000000000074696d65;
mem[142]<=80'h00000000000000006973;
mem[143]<=80'h0000000000000000003f;

//12th Sentence
mem[144]<=80'h0000000000004e657874;
mem[145]<=80'h00000000666c69676874;
mem[146]<=80'h0000000000000000746f;
mem[147]<=80'h00000000005065727468;
mem[148]<=80'h00000000000000006973;
mem[149]<=80'h00000000000000006174;
mem[150]<=80'h00000000000000000035;
mem[151]<=80'h0000000000000000706d;
mem[152]<=80'h0000000000000000002e;
mem[153]<=80'h00416c7465726e617465;
mem[154]<=80'h00000000666c69676874;
mem[155]<=80'h0000000000000000746f;
mem[156]<=80'h00000000005065727468;
mem[157]<=80'h0000000000000000003f;

//13th Sentence
mem[158]<=80'h00000000000043484452;
mem[159]<=80'h00000000000000006973;
mem[160]<=80'h0000006c6f6361746564;
mem[161]<=80'h00000000000000006174;
mem[162]<=80'h00000000000000004336;
mem[163]<=80'h0000000000000000002e;
mem[164]<=80'h00005265736561726368;
mem[165]<=80'h000000006f6666696365; 
mem[166]<=80'h00000000000000006973;
mem[167]<=80'h00000000000000006174;
mem[168]<=80'h0000000000000000003f;

//14th Sentence
mem[169]<=80'h00000000000000546865;
mem[170]<=80'h0000636f6d7075746572;
mem[171]<=80'h0000000000006e616d65;
mem[172]<=80'h00000000000000006973;
mem[173]<=80'h000000000000004d6178;
mem[174]<=80'h0000000000000000002e;
mem[175]<=80'h000000000000446f6573;
mem[176]<=80'h00000000000000746865;
mem[177]<=80'h0000636f6d7075746572;
mem[178]<=80'h00000000000068617665;
mem[179]<=80'h00000000000000000061;
mem[180]<=80'h0000000000006e616d65;
mem[181]<=80'h0000000000000000003f;

//15th Sentence
mem[182]<=80'h0000000000004e657874;
mem[183]<=80'h00000000457572656361;
mem[184]<=80'h636f6e666572656e6365;
mem[185]<=80'h00000068617070656e73;
mem[186]<=80'h0000000000000000696e;
mem[187]<=80'h00000000000032303139;
mem[188]<=80'h0000000000000000002e;
mem[189]<=80'h00000000436f6d696e67;
mem[190]<=80'h00000000457572656361;
mem[191]<=80'h636f6e666572656e6365;
mem[192]<=80'h00000068617070656e73;
mem[193]<=80'h0000000000000000696e;
mem[194]<=80'h0000000000000000003f;

//16th Sentence
mem[195]<=80'h00000000005468616e6b;
mem[196]<=80'h00000000000000796f75;
mem[197]<=80'h000065766572796f6e65;
mem[198]<=80'h0000000000000000002e;
mem[199]<=80'h0000436f6e636c756465;
mem[200]<=80'h00000000000000746865;
mem[201]<=80'h00000000006576656e74;
mem[202]<=80'h0000000000000000003f;

//17th Sentence
mem[203]<=80'h000000000000476f6f64;
mem[204]<=80'h0000006d6f726e696e67;
mem[205]<=80'h0000000000000000746f;
mem[206]<=80'h00000000000000616c6c;
mem[207]<=80'h0000000000000000002e;
mem[208]<=80'h00000000004772656574;
mem[209]<=80'h000065766572796f6e65;
mem[210]<=80'h00000000000000000021;

//18th Sentence
mem[211]<=80'h00000000000000000049;
mem[212]<=80'h0000000000000000616d;
mem[213]<=80'h00000000000066726f6d;
mem[214]<=80'h0000000000496e646961;
mem[215]<=80'h0000000000000000002e;
mem[216]<=80'h000000000000596f7572;
mem[217]<=80'h000000006e6174697665;
mem[218]<=80'h00000000000000006973;
mem[219]<=80'h00000000000000000021;

//19th Sentence
mem[220]<=80'h00000000000000000049;
mem[221]<=80'h0000000000000000616d;
mem[222]<=80'h00007374756479696e67;
mem[223]<=80'h00000000000000006174;
mem[224]<=80'h0000005461796c6f7273;
mem[225]<=80'h756e6976657273697479;
mem[226]<=80'h0000000000000000002e;
mem[227]<=80'h00000000005768696368;
mem[228]<=80'h756e6976657273697479;
mem[229]<=80'h00000000000000617265;
mem[230]<=80'h00000000000000796f75;
mem[231]<=80'h00007374756479696e67;
mem[232]<=80'h00000000000000006174;
mem[233]<=80'h00000000000000000021;

//20th Sentence
mem[234]<=80'h00000000000000596f75;
mem[235]<=80'h00000000000000617265;
mem[236]<=80'h00000077656c636f6d65;
mem[237]<=80'h0000000000000000002e;
mem[238]<=80'h00000000005468616e6b;
mem[239]<=80'h00000000000000796f75;
mem[240]<=80'h00000000000000666f72;
mem[241]<=80'h00000000000000746865;
mem[242]<=80'h00000064657461696c73;
mem[243]<=80'h0000000000000000003f;

//empty
mem[244]<=80'h00000000000000000020;
mem[245]<=80'h00000000000000000020;
mem[246]<=80'h00000000000000000020;
mem[247]<=80'h00000000000000000020;
mem[248]<=80'h00000000000000000020;
mem[249]<=80'h00000000000000000020;
mem[250]<=80'h00000000000000000020;
mem[251]<=80'h00000000000000000020;
mem[252]<=80'h00000000000000000020;
mem[253]<=80'h00000000000000000020;
mem[254]<=80'h00000000000000000020;
mem[255]<=80'h00000000000000000020;
end
else 
begin
mem[0]<=80'h00000000000000000020;
//1st Sentence
mem[1]<=80'h00000053616d73756e67;
mem[2]<=80'h00000000000000006973;
mem[3]<=80'h0000006c6f6361746564;
mem[4]<=80'h0000000000000000696e;
mem[5]<=80'h0000000000536f757468;
mem[6]<=80'h00000000004b6f726561;
mem[7]<=80'h0000000000000000002e;
mem[8]<=80'h00000000005768657265;
mem[9]<=80'h00000000000000006973;
mem[10]<=80'h00000053616d73756e67;
mem[11]<=80'h0000006c6f6361746564;
mem[12]<=80'h0000000000000000003f;
//2nd Sentence
mem[13]<=80'h000000000000004c6565;
mem[14]<=80'h00000000004279756e67;
mem[15]<=80'h00000000000000006973;
mem[16]<=80'h00000000000000746865;
mem[17]<=80'h000000666f756e646572;
mem[18]<=80'h00000000000000006f66;
mem[19]<=80'h00000053616d73756e67;
mem[20]<=80'h0000000000000000002e;
mem[21]<=80'h0000000000000057686f;
mem[22]<=80'h00000000000000006973;
mem[23]<=80'h00000000000000746865;
mem[24]<=80'h000000666f756e646572;
mem[25]<=80'h00000000000000006f66;
mem[26]<=80'h00000053616d73756e67;
mem[27]<=80'h0000000000000000003f;
//3rd Sentence
mem[28]<=80'h00000000000000546865;
mem[29]<=80'h00000063757272656e74;
mem[30]<=80'h0000000000666f637573;
mem[31]<=80'h00000000000000006f66;
mem[32]<=80'h00000053616d73756e67;
mem[33]<=80'h00000000000000006973;
mem[34]<=80'h0000000000536d617274;
mem[35]<=80'h0000000070686f6e6573;
mem[36]<=80'h0000000000000000002e;
mem[37]<=80'h00000000000057686174;
mem[38]<=80'h00000000000000006973;
mem[39]<=80'h00000000000000546865;
mem[40]<=80'h0000000000666f637573;
mem[41]<=80'h00000000000000006f66;
mem[42]<=80'h00000053616d73756e67;
mem[43]<=80'h0000000000000000003f;

//4th Sentence
mem[44]<=80'h00000000000000005336;
mem[45]<=80'h00000000000000776173;
mem[46]<=80'h000072656c6561736564;
mem[47]<=80'h0000000000000000696e;
mem[48]<=80'h00000000000032303135;
mem[49]<=80'h0000000000000000002e;
mem[50]<=80'h0000000000005768656e;
mem[51]<=80'h00000000000000776173;
mem[52]<=80'h00000000000000005336;
mem[53]<=80'h000072656c6561736564;
mem[54]<=80'h0000000000000000003f;

// 5th Sentence
mem[55]<=80'h00000000000000005336;
mem[56]<=80'h00000000000000686173;
mem[57]<=80'h000000416e64726f6964;
mem[58]<=80'h00000000000000004f53;
mem[59]<=80'h0000000000000000002e;
mem[60]<=80'h00000000005768696368;
mem[61]<=80'h00000000000000004f53;
mem[62]<=80'h00000000000000006973;
mem[63]<=80'h00000070726573656e74;
mem[64]<=80'h0000000000000000696e;
mem[65]<=80'h00000000000000005336;
mem[66]<=80'h0000000000000000003f;


//6th Sentence
mem[67]<=80'h00000053616d73756e67;
mem[68]<=80'h00000000000000006973;
mem[69]<=80'h00000000000000000061;
mem[70]<=80'h00000000676c6f62616c;
mem[71]<=80'h000000636f6d70616e79;
mem[72]<=80'h0000000000000000002e;
mem[73]<=80'h00000000000000004973;
mem[74]<=80'h00000053616d73756e67;
mem[75]<=80'h00000000000000000061;
mem[76]<=80'h00006e6174696f6e616c;
mem[77]<=80'h000000636f6d70616e79;
mem[78]<=80'h0000000000000000003f;

//7th Sentence
mem[79]<=80'h0000000000004d61696e;
mem[80]<=80'h636f6d70657469746f72;
mem[81]<=80'h00000000000000006f66;
mem[82]<=80'h00000053616d73756e67;
mem[83]<=80'h00000000000000006973;
mem[84]<=80'h00000000004170706c65;
mem[85]<=80'h0000000000000000002e;
mem[86]<=80'h00000000000000546865;
mem[87]<=80'h0000000000004d61696e;
mem[88]<=80'h636f6d70657469746f72;  
mem[89]<=80'h00000000000000006f66;   
mem[90]<=80'h00000053616d73756e67;
mem[91]<=80'h0000000000000000003f;

//8th Sentence
mem[92]<=80'h00000000000000005336;
mem[93]<=80'h0000000000636f737473;
mem[94]<=80'h00000000000031303030;
mem[95]<=80'h000052696e6767697473;
mem[96]<=80'h0000000000000000002e;
mem[97]<=80'h00000000000000486f77;
mem[98]<=80'h0000000000006d756368;
mem[99]<=80'h000000000000646f6573;
mem[100]<=80'h00000000000000005336;
mem[101]<=80'h000000000000636f7374;
mem[102]<=80'h0000000000000000003f;

//9th Sentence
mem[103]<=80'h00000000000000005336;
mem[104]<=80'h0000000000000052414d;
mem[105]<=80'h00000000000073697a65;
mem[106]<=80'h00000000000000006973;
mem[107]<=80'h00000000000000000033;
mem[108]<=80'h00000000000000004742;
mem[109]<=80'h0000000000000000002e;
mem[110]<=80'h00000000000054656c6c;
mem[111]<=80'h00000000000000746865;
mem[112]<=80'h0000000000000052414d;
mem[113]<=80'h00000000000073697a65;
mem[114]<=80'h00000000000000006f66;
mem[115]<=80'h00000000000000005336;
mem[116]<=80'h0000000000000000003f;

//10th Sentence
mem[117]<=80'h00000041697261736961;
mem[118]<=80'h0000000000006d61696e;
mem[119]<=80'h000000006f6666696365;
mem[120]<=80'h00000000000000006973;
mem[121]<=80'h0000006c6f6361746564;
mem[122]<=80'h0000000000000000696e;
mem[123]<=80'h00000000537562616e67;
mem[124]<=80'h0000000000004a617961;
mem[125]<=80'h0000000000000000002e;
mem[126]<=80'h00004169726173696173;
mem[127]<=80'h0000000000006d61696e;
mem[128]<=80'h000000006f6666696365;
mem[129]<=80'h00000000000000006973;
mem[130]<=80'h0000006c6f6361746564;
mem[131]<=80'h0000000000000000696e;
mem[132]<=80'h0000000000000000003f;

//11th Sentence
mem[133]<=80'h0000000000414b303231;
mem[134]<=80'h00000061727269766573;
mem[135]<=80'h0000000000000000696e;
mem[136]<=80'h00000000000000000034;
mem[137]<=80'h0000000000686f757273;
mem[138]<=80'h0000000000000000002e;
mem[139]<=80'h000000414b3032312773;
mem[140]<=80'h0000006172726976616c;
mem[141]<=80'h00000000000074696d65;
mem[142]<=80'h00000000000000006973;
mem[143]<=80'h0000000000000000003f;

//12th Sentence
mem[144]<=80'h0000000000004e657874;
mem[145]<=80'h00000000666c69676874;
mem[146]<=80'h0000000000000000746f;
mem[147]<=80'h00000000005065727468;
mem[148]<=80'h00000000000000006973;
mem[149]<=80'h00000000000000006174;
mem[150]<=80'h00000000000000000035;
mem[151]<=80'h0000000000000000706d;
mem[152]<=80'h0000000000000000002e;
mem[153]<=80'h00416c7465726e617465;
mem[154]<=80'h00000000666c69676874;
mem[155]<=80'h0000000000000000746f;
mem[156]<=80'h00000000005065727468;
mem[157]<=80'h0000000000000000003f;

//13th Sentence
mem[158]<=80'h00000000000043484452;
mem[159]<=80'h00000000000000006973;
mem[160]<=80'h0000006c6f6361746564;
mem[161]<=80'h00000000000000006174;
mem[162]<=80'h00000000000000004336;
mem[163]<=80'h0000000000000000002e;
mem[164]<=80'h00005265736561726368;
mem[165]<=80'h000000006f6666696365; 
mem[166]<=80'h00000000000000006973;
mem[167]<=80'h00000000000000006174;
mem[168]<=80'h0000000000000000003f;

//14th Sentence
mem[169]<=80'h00000000000000546865;
mem[170]<=80'h0000636f6d7075746572;
mem[171]<=80'h0000000000006e616d65;
mem[172]<=80'h00000000000000006973;
mem[173]<=80'h000000000000004d6178;
mem[174]<=80'h0000000000000000002e;
mem[175]<=80'h000000000000446f6573;
mem[176]<=80'h00000000000000746865;
mem[177]<=80'h0000636f6d7075746572;
mem[178]<=80'h00000000000068617665;
mem[179]<=80'h00000000000000000061;
mem[180]<=80'h0000000000006e616d65;
mem[181]<=80'h0000000000000000003f;

//15th Sentence
mem[182]<=80'h0000000000004e657874;
mem[183]<=80'h00000000457572656361;
mem[184]<=80'h636f6e666572656e6365;
mem[185]<=80'h00000068617070656e73;
mem[186]<=80'h0000000000000000696e;
mem[187]<=80'h00000000000032303139;
mem[188]<=80'h0000000000000000002e;
mem[189]<=80'h00000000436f6d696e67;
mem[190]<=80'h00000000457572656361;
mem[191]<=80'h636f6e666572656e6365;
mem[192]<=80'h00000068617070656e73;
mem[193]<=80'h0000000000000000696e;
mem[194]<=80'h0000000000000000003f;

//16th Sentence
mem[195]<=80'h00000000005468616e6b;
mem[196]<=80'h00000000000000796f75;
mem[197]<=80'h000065766572796f6e65;
mem[198]<=80'h0000000000000000002e;
mem[199]<=80'h0000436f6e636c756465;
mem[200]<=80'h00000000000000746865;
mem[201]<=80'h00000000006576656e74;
mem[202]<=80'h0000000000000000003f;

//17th Sentence
mem[203]<=80'h000000000000476f6f64;
mem[204]<=80'h0000006d6f726e696e67;
mem[205]<=80'h0000000000000000746f;
mem[206]<=80'h00000000000000616c6c;
mem[207]<=80'h0000000000000000002e;
mem[208]<=80'h00000000004772656574;
mem[209]<=80'h000065766572796f6e65;
mem[210]<=80'h00000000000000000021;

//18th Sentence
mem[211]<=80'h00000000000000000049;
mem[212]<=80'h0000000000000000616d;
mem[213]<=80'h00000000000066726f6d;
mem[214]<=80'h0000000000496e646961;
mem[215]<=80'h0000000000000000002e;
mem[216]<=80'h000000000000596f7572;
mem[217]<=80'h000000006e6174697665;
mem[218]<=80'h00000000000000006973;
mem[219]<=80'h00000000000000000021;

//19th Sentence
mem[220]<=80'h00000000000000000049;
mem[221]<=80'h0000000000000000616d;
mem[222]<=80'h00007374756479696e67;
mem[223]<=80'h00000000000000006174;
mem[224]<=80'h0000005461796c6f7273;
mem[225]<=80'h756e6976657273697479;
mem[226]<=80'h0000000000000000002e;
mem[227]<=80'h00000000005768696368;
mem[228]<=80'h756e6976657273697479;
mem[229]<=80'h00000000000000617265;
mem[230]<=80'h00000000000000796f75;
mem[231]<=80'h00007374756479696e67;
mem[232]<=80'h00000000000000006174;
mem[233]<=80'h00000000000000000021;

//20th Sentence
mem[234]<=80'h00000000000000596f75;
mem[235]<=80'h00000000000000617265;
mem[236]<=80'h00000077656c636f6d65;
mem[237]<=80'h0000000000000000002e;
mem[238]<=80'h00000000005468616e6b;
mem[239]<=80'h00000000000000796f75;
mem[240]<=80'h00000000000000666f72;
mem[241]<=80'h00000000000000746865;
mem[242]<=80'h00000064657461696c73;
mem[243]<=80'h0000000000000000003f;

//empty
mem[244]<=80'h00000000000000000020;
mem[245]<=80'h00000000000000000020;
mem[246]<=80'h00000000000000000020;
mem[247]<=80'h00000000000000000020;
mem[248]<=80'h00000000000000000020;
mem[249]<=80'h00000000000000000020;
mem[250]<=80'h00000000000000000020;
mem[251]<=80'h00000000000000000020;
mem[252]<=80'h00000000000000000020;
mem[253]<=80'h00000000000000000020;
mem[254]<=80'h00000000000000000020;
mem[255]<=80'h00000000000000000020;
out<=mem[address];
end
end
endmodule




























    

