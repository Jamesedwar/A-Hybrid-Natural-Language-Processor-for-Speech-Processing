module Qdict(clk, rst, out, val);
input          clk,rst;
input         [7:0]val; 
reg [79:0] mem [0:255];
output       [79:0]out;
reg           [2:0]cnt;
reg          [79:0]out;
wire         [7:0] add;
reg         [7:0] wadd;

assign add =(cnt==3'd0)? val:wadd;
always @(posedge clk or negedge rst)
begin
if (rst==0)
begin
cnt<=0;
wadd<=0;
end
else
begin
wadd<= add+8'd1;
cnt <= cnt+3'd1;
end
end


always @(posedge clk or negedge rst)
begin
if(rst==0)
begin
//1st Query
mem[0]<=80'h0000000000000000002e;
mem[1]<=80'h00000000005768657265;
mem[2]<=80'h00000000000000006973;
mem[3]<=80'h00000053616d73756e67;
mem[4]<=80'h0000006c6f6361746564;
mem[5]<=80'h0000000000000000003f;
mem[6]<=80'h00000000000000000020;
mem[7]<=80'h00000000000000000020;
//2nd Sentence
mem[8]<=80'h0000000000000000002e;
mem[9]<=80'h0000000000000057686f;
mem[10]<=80'h00000000000000006973;
mem[11]<=80'h00000000000000746865;
mem[12]<=80'h000000666f756e646572;
mem[13]<=80'h00000000000000006f66;
mem[14]<=80'h00000053616d73756e67;
mem[15]<=80'h0000000000000000003f;
//3rd Sentence
mem[16]<=80'h0000000000000000002e;
mem[17]<=80'h00000000000057686174;
mem[18]<=80'h00000000000000006973;
mem[19]<=80'h00000000000000546865;
mem[20]<=80'h0000000000666f637573;
mem[21]<=80'h00000000000000006f66;
mem[22]<=80'h00000053616d73756e67;
mem[23]<=80'h0000000000000000003f;
//4th Sentence
mem[24]<=80'h0000000000005768656e;
mem[25]<=80'h00000000000000776173;
mem[26]<=80'h00000000000000005336;
mem[27]<=80'h000072656c6561736564;
mem[28]<=80'h0000000000000000003f;
mem[29]<=80'h00000000000000000020;
mem[30]<=80'h00000000000000000020;
mem[31]<=80'h00000000000000000020;
// 5th Sentence
mem[32]<=80'h0000000000000000002e;
mem[33]<=80'h00000000005768696368;
mem[34]<=80'h00000000000000004f53;
mem[35]<=80'h00000000000000006973;
mem[36]<=80'h00000070726573656e74;
mem[37]<=80'h0000000000000000696e;
mem[38]<=80'h00000000000000005336;
mem[39]<=80'h0000000000000000003f;

//6th Sentence
mem[40]<=80'h0000000000000000002e;
mem[41]<=80'h00000000000000004973;
mem[42]<=80'h00000053616d73756e67;
mem[43]<=80'h00000000000000000061;
mem[44]<=80'h00006e6174696f6e616c;
mem[45]<=80'h000000636f6d70616e79;
mem[46]<=80'h0000000000000000003f;
mem[47]<=80'h00000000000000000020;
//7th Sentence
mem[48]<=80'h0000000000000000002e;
mem[49]<=80'h00000000000000546865;
mem[50]<=80'h0000000000004d61696e;
mem[51]<=80'h636f6d70657469746f72;  
mem[52]<=80'h00000000000000006f66;   
mem[53]<=80'h00000053616d73756e67;
mem[54]<=80'h0000000000000000003f;
mem[55]<=80'h00000000000000000020;
//8th Sentence
mem[56]<=80'h0000000000000000002e;
mem[57]<=80'h00000000000000486f77;
mem[58]<=80'h0000000000006d756368;
mem[59]<=80'h000000000000646f6573;
mem[60]<=80'h00000000000000005336;
mem[61]<=80'h000000000000636f7374;
mem[62]<=80'h0000000000000000003f;
mem[63]<=80'h00000000000000000020;
//9th Sentence
mem[64]<=80'h0000000000000000002e;
mem[65]<=80'h00000000000054656c6c;
mem[66]<=80'h00000000000000746865;
mem[67]<=80'h0000000000000052414d;
mem[68]<=80'h00000000000073697a65;
mem[69]<=80'h00000000000000006f66;
mem[70]<=80'h00000000000000005336;
mem[71]<=80'h0000000000000000003f;
//10th Sentence
mem[72]<=80'h0000000000000000002e;
mem[73]<=80'h00004169726173696173;
mem[74]<=80'h0000000000006d61696e;
mem[75]<=80'h000000006f6666696365;
mem[76]<=80'h00000000000000006973;
mem[77]<=80'h0000006c6f6361746564;
mem[78]<=80'h0000000000000000696e;
mem[79]<=80'h0000000000000000003f;

//11th Sentence
mem[80]<=80'h0000000000000000002e;
mem[81]<=80'h000000414b3032312773;
mem[82]<=80'h0000006172726976616c;
mem[83]<=80'h00000000000074696d65;
mem[84]<=80'h00000000000000006973;
mem[85]<=80'h0000000000000000003f;
mem[86]<=80'h00000000000000000020;
mem[87]<=80'h00000000000000000020;

//12th Sentence
mem[88]<=80'h0000000000000000002e;
mem[89]<=80'h00416c7465726e617465;
mem[90]<=80'h00000000666c69676874;
mem[91]<=80'h0000000000000000746f;
mem[92]<=80'h00000000005065727468;
mem[93]<=80'h0000000000000000003f;
mem[94]<=80'h00000000000000000020;
mem[95]<=80'h00000000000000000020;

//13th Sentence
mem[96]<=80'h0000000000000000002e;
mem[97]<=80'h00005265736561726368;
mem[98]<=80'h000000006f6666696365; 
mem[99]<=80'h00000000000000006973;
mem[100]<=80'h00000000000000006174;
mem[101]<=80'h0000000000000000003f;
mem[102]<=80'h00000000000000000020;
mem[103]<=80'h00000000000000000020;

//14th Sentence
mem[104]<=80'h0000000000000000002e;
mem[105]<=80'h000000000000446f6573;
mem[106]<=80'h00000000000000746865;
mem[107]<=80'h0000636f6d7075746572;
mem[108]<=80'h00000000000068617665;
mem[109]<=80'h00000000000000000061;
mem[110]<=80'h0000000000006e616d65;
mem[111]<=80'h0000000000000000003f;

//15th Sentence
mem[112]<=80'h0000000000000000002e;
mem[113]<=80'h00000000436f6d696e67;
mem[114]<=80'h00000000457572656361;
mem[115]<=80'h636f6e666572656e6365;
mem[116]<=80'h00000068617070656e73;
mem[117]<=80'h0000000000000000696e;
mem[118]<=80'h0000000000000000003f;
mem[119]<=80'h00000000000000000020;

//16th Sentence
mem[120]<=80'h0000000000000000002e;
mem[121]<=80'h0000436f6e636c756465;
mem[122]<=80'h00000000000000746865;
mem[123]<=80'h00000000006576656e74;
mem[124]<=80'h0000000000000000003f;
mem[125]<=80'h00000000000000000020;
mem[126]<=80'h00000000000000000020;
mem[127]<=80'h00000000000000000020;

//17th Sentence
mem[128]<=80'h0000000000000000002e;
mem[129]<=80'h00000000004772656574;
mem[130]<=80'h000065766572796f6e65;
mem[131]<=80'h0000000000000000003f;
mem[132]<=80'h00000000000000000020;
mem[133]<=80'h00000000000000000020;
mem[134]<=80'h00000000000000000020;
mem[135]<=80'h00000000000000000020;

//18th Sentence
mem[136]<=80'h0000000000000000002e;
mem[137]<=80'h000000000000596f7572;
mem[138]<=80'h000000006e6174697665;
mem[139]<=80'h00000000000000006973;
mem[140]<=80'h00000000000000000021;
mem[141]<=80'h00000000000000000020;
mem[142]<=80'h00000000000000000020;
mem[143]<=80'h00000000000000000020;

//19th Sentence
mem[144]<=80'h0000000000000000002e;
mem[145]<=80'h00000000005768696368;
mem[146]<=80'h756e6976657273697479;
mem[147]<=80'h00000000000000617265;
mem[148]<=80'h00000000000000796f75;
mem[149]<=80'h00000000000000006174;
mem[150]<=80'h00000000000000000021;
mem[151]<=80'h00000000000000000020;

//20th Sentence

mem[152]<=80'h0000000000000000002e;
mem[153]<=80'h00000000005468616e6b;
mem[154]<=80'h00000000000000796f75;
mem[155]<=80'h00000000000000666f72;
mem[156]<=80'h00000064657461696c73;
mem[157]<=80'h0000000000000000003f;
mem[158]<=80'h00000000000000000020;
mem[159]<=80'h00000000000000000020;
//empty
mem[160]<=80'h00000000000000000020;
mem[161]<=80'h00000000000000000020;
mem[162]<=80'h00000000000000000020;
mem[163]<=80'h00000000000000000020;
mem[164]<=80'h00000000000000000020;
mem[165]<=80'h00000000000000000020;
mem[166]<=80'h00000000000000000020;
mem[167]<=80'h00000000000000000020;
mem[168]<=80'h00000000000000000020;
mem[169]<=80'h00000000000000000020;
mem[170]<=80'h00000000000000000020;
mem[171]<=80'h00000000000000000020;
mem[172]<=80'h00000000000000000020;
mem[173]<=80'h00000000000000000020;
mem[174]<=80'h00000000000000000020;
mem[175]<=80'h00000000000000000020;
mem[176]<=80'h00000000000000000020;
mem[177]<=80'h00000000000000000020;
mem[178]<=80'h00000000000000000020;
mem[179]<=80'h00000000000000000020;
mem[180]<=80'h00000000000000000020;
mem[181]<=80'h00000000000000000020;
mem[182]<=80'h00000000000000000020;
mem[183]<=80'h00000000000000000020;
mem[184]<=80'h00000000000000000020;
mem[185]<=80'h00000000000000000020;
mem[186]<=80'h00000000000000000020;
mem[187]<=80'h00000000000000000020;
mem[188]<=80'h00000000000000000020;
mem[189]<=80'h00000000000000000020;
mem[190]<=80'h00000000000000000020;
mem[191]<=80'h00000000000000000020;
mem[192]<=80'h00000000000000000020;
mem[193]<=80'h00000000000000000020;
mem[194]<=80'h00000000000000000020;
mem[195]<=80'h00000000000000000020;
mem[196]<=80'h00000000000000000020;
mem[197]<=80'h00000000000000000020;
mem[198]<=80'h00000000000000000020;
mem[199]<=80'h00000000000000000020;
mem[200]<=80'h00000000000000000020;
mem[201]<=80'h00000000000000000020;
mem[202]<=80'h00000000000000000020;
mem[203]<=80'h00000000000000000020;
mem[204]<=80'h00000000000000000020;
mem[205]<=80'h00000000000000000020;
mem[206]<=80'h00000000000000000020;
mem[207]<=80'h00000000000000000020;
mem[208]<=80'h00000000000000000020;
mem[209]<=80'h00000000000000000020;
mem[210]<=80'h00000000000000000020;
mem[211]<=80'h00000000000000000020;
mem[212]<=80'h00000000000000000020;
mem[213]<=80'h00000000000000000020;
mem[214]<=80'h00000000000000000020;
mem[215]<=80'h00000000000000000020;
mem[216]<=80'h00000000000000000020;
mem[217]<=80'h00000000000000000020;
mem[218]<=80'h00000000000000000020;
mem[219]<=80'h00000000000000000020;
mem[220]<=80'h00000000000000000020;
mem[221]<=80'h00000000000000000020;
mem[222]<=80'h00000000000000000020;
mem[223]<=80'h00000000000000000020;
mem[224]<=80'h00000000000000000020;
mem[225]<=80'h00000000000000000020;
mem[226]<=80'h00000000000000000020;
mem[227]<=80'h00000000000000000020;
mem[228]<=80'h00000000000000000020;
mem[229]<=80'h00000000000000000020;
mem[230]<=80'h00000000000000000020;
mem[231]<=80'h00000000000000000020;
mem[232]<=80'h00000000000000000020;
mem[233]<=80'h00000000000000000020;
mem[234]<=80'h00000000000000000020;
mem[235]<=80'h00000000000000000020;
mem[236]<=80'h00000000000000000020;
mem[237]<=80'h00000000000000000020;
mem[238]<=80'h00000000000000000020;
mem[239]<=80'h00000000000000000020;
mem[240]<=80'h00000000000000000020;
mem[241]<=80'h00000000000000000020;
mem[242]<=80'h00000000000000000020;
mem[243]<=80'h00000000000000000020;
mem[244]<=80'h00000000000000000020;
mem[245]<=80'h00000000000000000020;
mem[246]<=80'h00000000000000000020;
mem[247]<=80'h00000000000000000020;
mem[248]<=80'h00000000000000000020;
mem[249]<=80'h00000000000000000020;
mem[250]<=80'h00000000000000000020;
mem[251]<=80'h00000000000000000020;
mem[252]<=80'h00000000000000000020;
mem[253]<=80'h00000000000000000020;
mem[254]<=80'h00000000000000000020;
mem[255]<=80'h00000000000000000020;
out<=0;
end
else
begin
//1st Query
mem[0]<=80'h0000000000000000002e;
mem[1]<=80'h00000000005768657265;
mem[2]<=80'h00000000000000006973;
mem[3]<=80'h00000053616d73756e67;
mem[4]<=80'h0000006c6f6361746564;
mem[5]<=80'h0000000000000000003f;
mem[6]<=80'h00000000000000000020;
mem[7]<=80'h00000000000000000020;
//2nd Sentence
mem[8]<=80'h0000000000000000002e;
mem[9]<=80'h0000000000000057686f;
mem[10]<=80'h00000000000000006973;
mem[11]<=80'h00000000000000746865;
mem[12]<=80'h000000666f756e646572;
mem[13]<=80'h00000000000000006f66;
mem[14]<=80'h00000053616d73756e67;
mem[15]<=80'h0000000000000000003f;
//3rd Sentence
mem[16]<=80'h0000000000000000002e;
mem[17]<=80'h00000000000057686174;
mem[18]<=80'h00000000000000006973;
mem[19]<=80'h00000000000000546865;
mem[20]<=80'h0000000000666f637573;
mem[21]<=80'h00000000000000006f66;
mem[22]<=80'h00000053616d73756e67;
mem[23]<=80'h0000000000000000003f;
//4th Sentence
mem[24]<=80'h0000000000005768656e;
mem[25]<=80'h00000000000000776173;
mem[26]<=80'h00000000000000005336;
mem[27]<=80'h000072656c6561736564;
mem[28]<=80'h0000000000000000003f;
mem[29]<=80'h00000000000000000020;
mem[30]<=80'h00000000000000000020;
mem[31]<=80'h00000000000000000020;
// 5th Sentence
mem[32]<=80'h0000000000000000002e;
mem[33]<=80'h00000000005768696368;
mem[34]<=80'h00000000000000004f53;
mem[35]<=80'h00000000000000006973;
mem[36]<=80'h00000070726573656e74;
mem[37]<=80'h0000000000000000696e;
mem[38]<=80'h00000000000000005336;
mem[39]<=80'h0000000000000000003f;

//6th Sentence
mem[40]<=80'h0000000000000000002e;
mem[41]<=80'h00000000000000004973;
mem[42]<=80'h00000053616d73756e67;
mem[43]<=80'h00000000000000000061;
mem[44]<=80'h00006e6174696f6e616c;
mem[45]<=80'h000000636f6d70616e79;
mem[46]<=80'h0000000000000000003f;
mem[47]<=80'h00000000000000000020;
//7th Sentence
mem[48]<=80'h0000000000000000002e;
mem[49]<=80'h00000000000000546865;
mem[50]<=80'h0000000000004d61696e;
mem[51]<=80'h636f6d70657469746f72;  
mem[52]<=80'h00000000000000006f66;   
mem[53]<=80'h00000053616d73756e67;
mem[54]<=80'h0000000000000000003f;
mem[55]<=80'h00000000000000000020;
//8th Sentence
mem[56]<=80'h0000000000000000002e;
mem[57]<=80'h00000000000000486f77;
mem[58]<=80'h0000000000006d756368;
mem[59]<=80'h000000000000646f6573;
mem[60]<=80'h00000000000000005336;
mem[61]<=80'h000000000000636f7374;
mem[62]<=80'h0000000000000000003f;
mem[63]<=80'h00000000000000000020;
//9th Sentence
mem[64]<=80'h0000000000000000002e;
mem[65]<=80'h00000000000054656c6c;
mem[66]<=80'h00000000000000746865;
mem[67]<=80'h0000000000000052414d;
mem[68]<=80'h00000000000073697a65;
mem[69]<=80'h00000000000000006f66;
mem[70]<=80'h00000000000000005336;
mem[71]<=80'h0000000000000000003f;
//10th Sentence
mem[72]<=80'h0000000000000000002e;
mem[73]<=80'h00004169726173696173;
mem[74]<=80'h0000000000006d61696e;
mem[75]<=80'h000000006f6666696365;
mem[76]<=80'h00000000000000006973;
mem[77]<=80'h0000006c6f6361746564;
mem[78]<=80'h0000000000000000696e;
mem[79]<=80'h0000000000000000003f;

//11th Sentence
mem[80]<=80'h0000000000000000002e;
mem[81]<=80'h000000414b3032312773;
mem[82]<=80'h0000006172726976616c;
mem[83]<=80'h00000000000074696d65;
mem[84]<=80'h00000000000000006973;
mem[85]<=80'h0000000000000000003f;
mem[86]<=80'h00000000000000000020;
mem[87]<=80'h00000000000000000020;

//12th Sentence
mem[88]<=80'h0000000000000000002e;
mem[89]<=80'h00416c7465726e617465;
mem[90]<=80'h00000000666c69676874;
mem[91]<=80'h0000000000000000746f;
mem[92]<=80'h00000000005065727468;
mem[93]<=80'h0000000000000000003f;
mem[94]<=80'h00000000000000000020;
mem[95]<=80'h00000000000000000020;

//13th Sentence
mem[96]<=80'h0000000000000000002e;
mem[97]<=80'h00005265736561726368;
mem[98]<=80'h000000006f6666696365; 
mem[99]<=80'h00000000000000006973;
mem[100]<=80'h00000000000000006174;
mem[101]<=80'h0000000000000000003f;
mem[102]<=80'h00000000000000000020;
mem[103]<=80'h00000000000000000020;

//14th Sentence
mem[104]<=80'h0000000000000000002e;
mem[105]<=80'h000000000000446f6573;
mem[106]<=80'h00000000000000746865;
mem[107]<=80'h0000636f6d7075746572;
mem[108]<=80'h00000000000068617665;
mem[109]<=80'h00000000000000000061;
mem[110]<=80'h0000000000006e616d65;
mem[111]<=80'h0000000000000000003f;

//15th Sentence
mem[112]<=80'h0000000000000000002e;
mem[113]<=80'h00000000436f6d696e67;
mem[114]<=80'h00000000457572656361;
mem[115]<=80'h636f6e666572656e6365;
mem[116]<=80'h00000068617070656e73;
mem[117]<=80'h0000000000000000696e;
mem[118]<=80'h0000000000000000003f;
mem[119]<=80'h00000000000000000020;

//16th Sentence
mem[120]<=80'h0000000000000000002e;
mem[121]<=80'h0000436f6e636c756465;
mem[122]<=80'h00000000000000746865;
mem[123]<=80'h00000000006576656e74;
mem[124]<=80'h0000000000000000003f;
mem[125]<=80'h00000000000000000020;
mem[126]<=80'h00000000000000000020;
mem[127]<=80'h00000000000000000020;

//17th Sentence
mem[128]<=80'h0000000000000000002e;
mem[129]<=80'h00000000004772656574;
mem[130]<=80'h000065766572796f6e65;
mem[131]<=80'h0000000000000000003f;
mem[132]<=80'h00000000000000000020;
mem[133]<=80'h00000000000000000020;
mem[134]<=80'h00000000000000000020;
mem[135]<=80'h00000000000000000020;

//18th Sentence
mem[136]<=80'h0000000000000000002e;
mem[137]<=80'h000000000000596f7572;
mem[138]<=80'h000000006e6174697665;
mem[139]<=80'h00000000000000006973;
mem[140]<=80'h00000000000000000021;
mem[141]<=80'h00000000000000000020;
mem[142]<=80'h00000000000000000020;
mem[143]<=80'h00000000000000000020;

//19th Sentence
mem[144]<=80'h0000000000000000002e;
mem[145]<=80'h00000000005768696368;
mem[146]<=80'h756e6976657273697479;
mem[147]<=80'h00000000000000617265;
mem[148]<=80'h00000000000000796f75;
mem[149]<=80'h00000000000000006174;
mem[150]<=80'h00000000000000000021;
mem[151]<=80'h00000000000000000020;

//20th Sentence

mem[152]<=80'h0000000000000000002e;
mem[153]<=80'h00000000005468616e6b;
mem[154]<=80'h00000000000000796f75;
mem[155]<=80'h00000000000000666f72;
mem[156]<=80'h00000064657461696c73;
mem[157]<=80'h0000000000000000003f;
mem[158]<=80'h00000000000000000020;
mem[159]<=80'h00000000000000000020;
//empty
mem[160]<=80'h00000000000000000020;
mem[161]<=80'h00000000000000000020;
mem[162]<=80'h00000000000000000020;
mem[163]<=80'h00000000000000000020;
mem[164]<=80'h00000000000000000020;
mem[165]<=80'h00000000000000000020;
mem[166]<=80'h00000000000000000020;
mem[167]<=80'h00000000000000000020;
mem[168]<=80'h00000000000000000020;
mem[169]<=80'h00000000000000000020;
mem[170]<=80'h00000000000000000020;
mem[171]<=80'h00000000000000000020;
mem[172]<=80'h00000000000000000020;
mem[173]<=80'h00000000000000000020;
mem[174]<=80'h00000000000000000020;
mem[175]<=80'h00000000000000000020;
mem[176]<=80'h00000000000000000020;
mem[177]<=80'h00000000000000000020;
mem[178]<=80'h00000000000000000020;
mem[179]<=80'h00000000000000000020;
mem[180]<=80'h00000000000000000020;
mem[181]<=80'h00000000000000000020;
mem[182]<=80'h00000000000000000020;
mem[183]<=80'h00000000000000000020;
mem[184]<=80'h00000000000000000020;
mem[185]<=80'h00000000000000000020;
mem[186]<=80'h00000000000000000020;
mem[187]<=80'h00000000000000000020;
mem[188]<=80'h00000000000000000020;
mem[189]<=80'h00000000000000000020;
mem[190]<=80'h00000000000000000020;
mem[191]<=80'h00000000000000000020;
mem[192]<=80'h00000000000000000020;
mem[193]<=80'h00000000000000000020;
mem[194]<=80'h00000000000000000020;
mem[195]<=80'h00000000000000000020;
mem[196]<=80'h00000000000000000020;
mem[197]<=80'h00000000000000000020;
mem[198]<=80'h00000000000000000020;
mem[199]<=80'h00000000000000000020;
mem[200]<=80'h00000000000000000020;
mem[201]<=80'h00000000000000000020;
mem[202]<=80'h00000000000000000020;
mem[203]<=80'h00000000000000000020;
mem[204]<=80'h00000000000000000020;
mem[205]<=80'h00000000000000000020;
mem[206]<=80'h00000000000000000020;
mem[207]<=80'h00000000000000000020;
mem[208]<=80'h00000000000000000020;
mem[209]<=80'h00000000000000000020;
mem[210]<=80'h00000000000000000020;
mem[211]<=80'h00000000000000000020;
mem[212]<=80'h00000000000000000020;
mem[213]<=80'h00000000000000000020;
mem[214]<=80'h00000000000000000020;
mem[215]<=80'h00000000000000000020;
mem[216]<=80'h00000000000000000020;
mem[217]<=80'h00000000000000000020;
mem[218]<=80'h00000000000000000020;
mem[219]<=80'h00000000000000000020;
mem[220]<=80'h00000000000000000020;
mem[221]<=80'h00000000000000000020;
mem[222]<=80'h00000000000000000020;
mem[223]<=80'h00000000000000000020;
mem[224]<=80'h00000000000000000020;
mem[225]<=80'h00000000000000000020;
mem[226]<=80'h00000000000000000020;
mem[227]<=80'h00000000000000000020;
mem[228]<=80'h00000000000000000020;
mem[229]<=80'h00000000000000000020;
mem[230]<=80'h00000000000000000020;
mem[231]<=80'h00000000000000000020;
mem[232]<=80'h00000000000000000020;
mem[233]<=80'h00000000000000000020;
mem[234]<=80'h00000000000000000020;
mem[235]<=80'h00000000000000000020;
mem[236]<=80'h00000000000000000020;
mem[237]<=80'h00000000000000000020;
mem[238]<=80'h00000000000000000020;
mem[239]<=80'h00000000000000000020;
mem[240]<=80'h00000000000000000020;
mem[241]<=80'h00000000000000000020;
mem[242]<=80'h00000000000000000020;
mem[243]<=80'h00000000000000000020;
mem[244]<=80'h00000000000000000020;
mem[245]<=80'h00000000000000000020;
mem[246]<=80'h00000000000000000020;
mem[247]<=80'h00000000000000000020;
mem[248]<=80'h00000000000000000020;
mem[249]<=80'h00000000000000000020;
mem[250]<=80'h00000000000000000020;
mem[251]<=80'h00000000000000000020;
mem[252]<=80'h00000000000000000020;
mem[253]<=80'h00000000000000000020;
mem[254]<=80'h00000000000000000020;
mem[255]<=80'h00000000000000000020;
out <=  mem[wadd];
end
end
endmodule