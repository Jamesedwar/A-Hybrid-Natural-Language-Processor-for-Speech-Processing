module SigmoidROM(out, add, CS, read); 
output[7:0] out;
input[7:0] add;
input CS,read;
reg [7:0] out;
reg [7:0] ROM[0:255];
always @(posedge CS)
begin
ROM[0] <= 8'd255;	
ROM[1] <= 8'd254;
ROM[2] <= 8'd253; 
ROM[3] <= 8'd252;
ROM[4] <= 8'd251;
ROM[5] <= 8'd250;
ROM[6] <= 8'd249;
ROM[7] <= 8'd248;
ROM[8] <= 8'd247;
ROM[9] <= 8'd246;
ROM[10] <= 8'd245;
ROM[11] <= 8'd244;
ROM[12] <= 8'd243;
ROM[13] <= 8'd242;
ROM[14] <= 8'd241;
ROM[15] <= 8'd240;
ROM[16] <= 8'd239;
ROM[17] <= 8'd238;
ROM[18] <= 8'd237;
ROM[19] <= 8'd236;
ROM[20] <= 8'd235;
ROM[21] <= 8'd234;
ROM[22] <= 8'd233;
ROM[23] <= 8'd232;
ROM[24] <= 8'd231;
ROM[25] <= 8'd230;
ROM[26] <= 8'd229;
ROM[27] <= 8'd228;
ROM[28] <= 8'd227;
ROM[29] <= 8'd226;
ROM[30] <= 8'd225;
ROM[31] <= 8'd224;
ROM[32] <= 8'd223;
ROM[33] <= 8'd222;
ROM[34] <= 8'd221;
ROM[35] <= 8'd220;
ROM[36] <= 8'd219;
ROM[37] <= 8'd218;
ROM[38] <= 8'd217;
ROM[39] <= 8'd216;
ROM[40] <= 8'd215;
ROM[41] <= 8'd214;
ROM[42] <= 8'd213;
ROM[43] <= 8'd212;
ROM[44] <= 8'd211;
ROM[45] <= 8'd210;
ROM[46] <= 8'd209;
ROM[47] <= 8'd208;
ROM[48] <= 8'd207;
ROM[49] <= 8'd206;
ROM[50] <= 8'd205;
ROM[51] <= 8'd204;
ROM[52] <= 8'd203;
ROM[53] <= 8'd202;
ROM[54] <= 8'd201;
ROM[55] <= 8'd200;
ROM[56] <= 8'd199;
ROM[57] <= 8'd198;
ROM[58] <= 8'd197;
ROM[59] <= 8'd196;
ROM[60] <= 8'd195;
ROM[61] <= 8'd194;
ROM[62] <= 8'd193;
ROM[63] <= 8'd192;
ROM[64] <= 8'd191;
ROM[65] <= 8'd190;
ROM[66] <= 8'd189;
ROM[67] <= 8'd188;
ROM[68] <= 8'd187;
ROM[69] <= 8'd186;
ROM[70] <= 8'd185;
ROM[71] <= 8'd184;
ROM[72] <= 8'd183;
ROM[73] <= 8'd182;
ROM[74] <= 8'd181;
ROM[75] <= 8'd180;
ROM[76] <= 8'd179;
ROM[77] <= 8'd178;
ROM[78] <= 8'd177;
ROM[79] <= 8'd176;
ROM[80] <= 8'd175;
ROM[81] <= 8'd174;
ROM[82] <= 8'd173;
ROM[83] <= 8'd172;
ROM[84] <= 8'd171;
ROM[85] <= 8'd170;
ROM[86] <= 8'd169;
ROM[87] <= 8'd168;
ROM[88] <= 8'd167;
ROM[89] <= 8'd166;
ROM[90] <= 8'd165;
ROM[91] <= 8'd164;
ROM[92] <= 8'd163;
ROM[93] <= 8'd162;
ROM[94] <= 8'd161;
ROM[95] <= 8'd160;
ROM[96] <= 8'd159;
ROM[97] <= 8'd158;
ROM[98] <= 8'd157;			
ROM[99] <= 8'd156;
ROM[100] <= 8'd155;
ROM[101] <= 8'd154;
ROM[102] <= 8'd153;
ROM[103] <= 8'd152;
ROM[104] <= 8'd151;
ROM[105] <= 8'd150;
ROM[106] <= 8'd149;
ROM[107] <= 8'd148;
ROM[108] <= 8'd147;	
ROM[109] <= 8'd146;
ROM[110] <= 8'd145;
ROM[111] <= 8'd144;
ROM[112] <= 8'd143;
ROM[113] <= 8'd142;
ROM[114] <= 8'd141;
ROM[115] <= 8'd140;
ROM[116] <= 8'd139;
ROM[117] <= 8'd138;
ROM[118] <= 8'd137;
ROM[119] <= 8'd136;
ROM[120] <= 8'd135;
ROM[121] <= 8'd134;
ROM[122] <= 8'd133;
ROM[123] <= 8'd132;
ROM[124] <= 8'd131;
ROM[125] <= 8'd130;
ROM[126] <= 8'd129;
ROM[127] <= 8'd128;	
ROM[128] <= 8'd127;
ROM[129] <= 8'd126; 
ROM[130] <= 8'd125;
ROM[131] <= 8'd124;
ROM[132] <= 8'd123;
ROM[133] <= 8'd122;
ROM[134] <= 8'd121;
ROM[135] <= 8'd120;
ROM[136] <= 8'd119;
ROM[137] <= 8'd118;
ROM[138] <= 8'd117;
ROM[139] <= 8'd116;
ROM[140] <= 8'd115;
ROM[141] <= 8'd114;
ROM[142] <= 8'd113;
ROM[143] <= 8'd112;
ROM[144] <= 8'd111;
ROM[145] <= 8'd110;
ROM[146] <= 8'd109;
ROM[147] <= 8'd108;
ROM[148] <= 8'd107;
ROM[149] <= 8'd106;
ROM[150] <= 8'd105;
ROM[151] <= 8'd104;
ROM[152] <= 8'd103;
ROM[153] <= 8'd102;
ROM[154] <= 8'd101;
ROM[155] <= 8'd100;
ROM[156] <= 8'd99;
ROM[157] <= 8'd98;
ROM[158] <= 8'd97;
ROM[159] <= 8'd96;
ROM[160] <= 8'd95;
ROM[161] <= 8'd94;
ROM[162] <= 8'd93;
ROM[163] <= 8'd92;
ROM[164] <= 8'd91;
ROM[165] <= 8'd90;
ROM[166] <= 8'd89;
ROM[167] <= 8'd88;
ROM[168] <= 8'd87;
ROM[169] <= 8'd86;
ROM[170] <= 8'd85;
ROM[171] <= 8'd84;
ROM[172] <= 8'd83;
ROM[173] <= 8'd82;
ROM[174] <= 8'd81;
ROM[175] <= 8'd80;
ROM[176] <= 8'd79;
ROM[177] <= 8'd78;
ROM[178] <= 8'd77;
ROM[179] <= 8'd76;
ROM[180] <= 8'd75;
ROM[181] <= 8'd74;
ROM[182] <= 8'd73;
ROM[183] <= 8'd72;
ROM[184] <= 8'd71;
ROM[185] <= 8'd70;
ROM[186] <= 8'd69;
ROM[187] <= 8'd68;
ROM[188] <= 8'd67;
ROM[189] <= 8'd66;
ROM[190] <= 8'd65;
ROM[191] <= 8'd64;
ROM[192] <= 8'd63;
ROM[193] <= 8'd62;
ROM[194] <= 8'd61;
ROM[195] <= 8'd60;
ROM[196] <= 8'd59;
ROM[197] <= 8'd58;
ROM[198] <= 8'd57;
ROM[199] <= 8'd56;
ROM[200] <= 8'd55;
ROM[201] <= 8'd54;
ROM[202] <= 8'd53;
ROM[203] <= 8'd52;
ROM[204] <= 8'd51;
ROM[205] <= 8'd50;
ROM[206] <= 8'd49;
ROM[207] <= 8'd48;
ROM[208] <= 8'd47;
ROM[209] <= 8'd46;
ROM[210] <= 8'd45;
ROM[211] <= 8'd44;
ROM[212] <= 8'd43;
ROM[213] <= 8'd42;
ROM[214] <= 8'd41;
ROM[215] <= 8'd40;
ROM[216] <= 8'd39;
ROM[217] <= 8'd38;
ROM[218] <= 8'd37;
ROM[219] <= 8'd36;
ROM[220] <= 8'd35;
ROM[221] <= 8'd34;
ROM[222] <= 8'd33;
ROM[223] <= 8'd32;
ROM[224] <= 8'd31;
ROM[225] <= 8'd30;			
ROM[226] <= 8'd29;
ROM[227] <= 8'd28;
ROM[228] <= 8'd27;
ROM[229] <= 8'd26;
ROM[230] <= 8'd25;
ROM[231] <= 8'd24;
ROM[232] <= 8'd23;
ROM[233] <= 8'd22;
ROM[234] <= 8'd21;
ROM[235] <= 8'd20;	
ROM[236] <= 8'd19;
ROM[237] <= 8'd18;
ROM[238] <= 8'd17;
ROM[239] <= 8'd16;
ROM[240] <= 8'd15;
ROM[241] <= 8'd14;
ROM[242] <= 8'd13;
ROM[243] <= 8'd12;
ROM[244] <= 8'd11;
ROM[245] <= 8'd10;
ROM[246] <= 8'd09;
ROM[247] <= 8'd08;
ROM[248] <= 8'd07;
ROM[249] <= 8'd06;
ROM[250] <= 8'd05;
ROM[251] <= 8'd04;
ROM[252] <= 8'd03;
ROM[253] <= 8'd02;
ROM[254] <= 8'd01;
ROM[255] <= 8'd00;
if(read==1)
out<=ROM[add];
else 
out<=0;
end
endmodule