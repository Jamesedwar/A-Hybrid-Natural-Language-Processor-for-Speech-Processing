module Hexa_Key_Encoder(in, out, en);
input en;

input [79:0]in;
output [7:0]out;


reg[7:0]out;
always@(en or in)
begin
if(en==0)
out<=0;
else
begin
case(in)
80'h00000000000000000020:out<=8'd0;
80'h00000053616d73756e67:out<=8'd1;
80'h00000000000000006973:out<=8'd2;
80'h0000006c6f6361746564:out<=8'd3;
80'h0000000000000000696e:out<=8'd4;
80'h0000000000536f757468:out<=8'd5;
80'h00000000004b6f726561:out<=8'd6;
80'h0000000000000000002e:out<=8'd7;
80'h00000000005768657265:out<=8'd8;
80'h0000000000000000003f:out<=8'd9;
80'h000000000000004c6565:out<=8'd10;
80'h00000000004279756e67:out<=8'd11;
80'h00000000000000746865:out<=8'd12;
80'h000000666f756e646572:out<=8'd13;
80'h00000000000000006f66:out<=8'd14;
80'h00000000000000546865:out<=8'd15;
80'h0000000000000057686f:out<=8'd16;
80'h00000063757272656e74:out<=8'd17;
80'h0000000000666f637573:out<=8'd18;
80'h0000000000536d617274:out<=8'd19;
80'h0000000070686f6e6573:out<=8'd20;
80'h00000000000057686174:out<=8'd21;
80'h00000000000000005336:out<=8'd22;
80'h00000000000000776173:out<=8'd23;
80'h000072656c6561736564:out<=8'd24;
80'h00000000000032303135:out<=8'd25;
80'h0000000000005768656e:out<=8'd26;
80'h00000000000000686173:out<=8'd27;
80'h000000416e64726f6964:out<=8'd28;
80'h00000000000000004f53:out<=8'd29;
80'h00000000005768696368:out<=8'd30;
80'h00000070726573656e74:out<=8'd31;
80'h00000000000000000061:out<=8'd32;
80'h00000000676c6f62616c:out<=8'd33;
80'h000000636f6d70616e79:out<=8'd34;
80'h00000000000000004973:out<=8'd35;
80'h00006e6174696f6e616c:out<=8'd36;
80'h0000000000004d61696e:out<=8'd37;
80'h636f6d70657469746f72:out<=8'd38;
80'h00000000004170706c65:out<=8'd39;
80'h0000000000636f737473:out<=8'd40;
80'h00000000000031303030:out<=8'd41;
80'h000052696e6767697473:out<=8'd42;
80'h00000000000000486f77:out<=8'd43;
80'h0000000000006d756368:out<=8'd44;
80'h000000000000646f6573:out<=8'd45;
80'h000000000000636f7374:out<=8'd46;
80'h0000000000000052414d:out<=8'd47;
80'h00000000000073697a65:out<=8'd48;
80'h00000000000000000033:out<=8'd49;
80'h00000000000000004742:out<=8'd50;
80'h00000000000054656c6c:out<=8'd51;
80'h00000041697261736961:out<=8'd52;
80'h0000000000006d61696e:out<=8'd53;
80'h000000006f6666696365:out<=8'd54;
80'h00000000537562616e67:out<=8'd55;
80'h0000000000004a617961:out<=8'd56;
80'h00416972617369612773:out<=8'd57;
80'h0000000000414b303231:out<=8'd58;
80'h00000061727269766573:out<=8'd59;
80'h00000000000000000034:out<=8'd60;
80'h0000000000686f757273:out<=8'd61;
80'h000000414b3032312773:out<=8'd62;
80'h0000006172726976616c:out<=8'd63;
80'h00000000000074696d65:out<=8'd64;
80'h0000000000004e657874:out<=8'd65;
80'h00000000000072756e73:out<=8'd66;
80'h00000000666c69676874:out<=8'd67;
80'h00000000005065727468:out<=8'd68;
80'h00000000000000006174:out<=8'd69;
80'h00000000000000000035:out<=8'd70;
80'h0000000000000000706d:out<=8'd71;
80'h00416c7465726e617465:out<=8'd72;
80'h00000000000043484452:out<=8'd73;
80'h00000000000000004336:out<=8'd74;
80'h00005265736561726368:out<=8'd75;
80'h0000000000006e616d65:out<=8'd76;
80'h000000000000004d6178:out<=8'd77;
80'h000000000000446f6573:out<=8'd78;
80'h00000000000068617665:out<=8'd79;
80'h00000000457572656361:out<=8'd80;
80'h636f6e666572656e6365:out<=8'd81;
80'h00000068617070656e73:out<=8'd82;
80'h00000000000032303139:out<=8'd83;
80'h00000000436f6d696e67:out<=8'd84;
80'h00000000005468616e6b:out<=8'd85;
80'h00000000000000796f75:out<=8'd86;
80'h000065766572796f6e65:out<=8'd87;
80'h0000436f6e636c756465:out<=8'd88;
80'h00000000006576656e74:out<=8'd89;
80'h000000000000476f6f64:out<=8'd90;
80'h0000006d6f726e696e67:out<=8'd91;
80'h00000000000000616c6c:out<=8'd92;
80'h00000000004772656574:out<=8'd93;
80'h0000000000000000616d:out<=8'd94;
80'h00000000000066726f6d:out<=8'd95;
80'h0000000000496e646961:out<=8'd96;
80'h000000000000596f7572:out<=8'd97;
80'h000000006e6174697665:out<=8'd98;
80'h00007374756479696e67:out<=8'd99;
80'h0000005461796c6f7273:out<=8'd100;
80'h756e6976657273697479:out<=8'd101;
80'h00000000000000617265:out<=8'd102;
80'h00000077656c636f6d65:out<=8'd103;

default:out<=8'd00;
endcase
end
end
endmodule
























    

